module EX_MEM_FF(, clk, rst_n, stall);

endmodule