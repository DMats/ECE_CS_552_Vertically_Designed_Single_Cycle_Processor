module ID();

endmodule
