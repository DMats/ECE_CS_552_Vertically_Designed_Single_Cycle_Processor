// Hazard Detect Module
// Author:  David Mateo
// This module is meant to contain all modules relating to hazard
// detect and control logic.
module HD(instr);

endmodule